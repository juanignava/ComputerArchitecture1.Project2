module alu_tb ();
	
	logic clk;
	logic [31:0] A, B;
	logic [2:0] sel;
	logic [31:0] C;
	logic flagZ;
	
	alu alu_TB (A, B, sel, C, flagZ);
	
	initial begin
		
		clk = 0; #2;
		
		// Suma, test 1:
		A = 32'b00000000000000000000000000000100; 
		B = 32'b00000000000000000000000000000011; sel = 3'b000; #2
		
		// Resta, test 1:
		A = 32'b00000000000000000000000000000100; 
		B = 32'b00000000000000000000000000000011; sel = 3'b001; #2
		
		// Multiplicación, test 1:
		A = 32'b00000000000000000000000000000100; 
		B = 32'b00000000000000000000000000000011; sel = 3'b010; #2
		
		// División entera, test 1:
		A = 32'b00000000000000000000000000000100; 
		B = 32'b00000000000000000000000000000011; sel = 3'b011; #2
		
		// División entera, test 2:
		A = 32'b00000000000000000000000000001000; 
		B = 32'b00000000000000000000000000000011; sel = 3'b011; #2
		
		// División entera, test 3:
		A = 32'b00000000000000000000000000101101; 
		B = 32'b00000000000000000000000000001001; sel = 3'b011; #2
		
		// Residuo, test 1:
		A = 32'b00000000000000000000000000000100; 
		B = 32'b00000000000000000000000000000011; sel = 3'b100; #2
		
		// Residuo, test 2:
		A = 32'b00000000000000000000000000001000; 
		B = 32'b00000000000000000000000000000011; sel = 3'b100; #2
		
		// Residuo, test 3:
		A = 32'b00000000000000000000000000101101; 
		B = 32'b00000000000000000000000000001001; sel = 3'b100; #2;
		
	end
	
	always begin
		clk=!clk; #1;
	end
	
endmodule